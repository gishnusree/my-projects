interface mux_if();
  logic [7:0] a, b, y;
  logic sel;
endinterface
